INFO:HDLCompiler:1061 - Parsing VHDL file "H:/zn/Projects/UV_Logger/readout/FPGA/uvl_readout/sources/com_dac_enc.vhd" into library work
INFO:ProjectMgmt - Parsing design hierarchy completed successfully.
INFO:HDLCompiler:1061 - Parsing VHDL file "H:/zn/Projects/UV_Logger/readout/FPGA/uvl_readout/sources/com_dac_enc.vhd" into library work
INFO:ProjectMgmt - Parsing design hierarchy completed successfully.
WARNING:ProjectMgmt - File H:/zn/Projects/UV_Logger/readout/FPGA/uvl_readout/uvl_readout_01_top.bit is missing.
